// $Id: $
// File name:   rcv_fifo_fsm.sv
// Created:     4/8/2017
// Author:      Natat Sombuntham
// Lab Section: 337-03
// Version:     1.0  Initial Design Entry
// Description: Implementation of rcv fifo fsm.
module rcv_fifo_fsm
(
	input wire clk,
	input wire n_rst,
	input wire rcv_enq_word,
	input wire full,
	input wire [1:0] tail_side,
	input wire fix_error,
	output reg count_en1,
	output reg sync_clr,
	output reg count_en2,
	output reg WE
);
//	typedef enum bit [2:0] {IDLE, WRITE, INC_IDX, INC_BOTH, FIX} stateType;
	typedef enum bit [1:0] {IDLE, INC_IDX, INC_BOTH, FIX} stateType;
	stateType state;
	stateType nextState;
	always_ff @ (negedge n_rst, posedge clk) begin : REG_LOGIC
		if (n_rst == 1'b0) begin
			state <= IDLE;
		end else begin
			state <= nextState;
		end
	end
	always_comb begin: NXT_LOGIC
		nextState = state;
		case (state)
			IDLE: begin
				if (rcv_enq_word && !full && tail_side != 3) begin
					nextState = INC_IDX;
				end
				else if (rcv_enq_word && !full && tail_side == 3) begin
					nextState = INC_BOTH;
				end
				else if (fix_error) begin
					nextState = FIX;
				end
			end
			INC_IDX: begin
				if (rcv_enq_word && !full && tail_side != 2) begin
					nextState = INC_IDX;
				end
				else if (rcv_enq_word && !full) begin
					nextState = INC_BOTH;
				end
				else begin
					nextState = IDLE;
				end
			end
			INC_BOTH: begin
				if (rcv_enq_word && !full) begin
					nextState = INC_IDX;
				end
				else begin
					nextState = IDLE;
				end
			end
			FIX: begin
				nextState = IDLE;
			end
		endcase
	end
	always_comb begin: OUTPUT_LOGIC
		count_en1 = 1'b0;
		sync_clr = 1'b0;
		count_en2 = 1'b0;
		WE = 1'b0;
		case (state)
			IDLE: begin
				//do nothing
			end
			INC_IDX: begin
				count_en1 = 1'b1;
				WE = 1'b1;
			end
			INC_BOTH: begin
				count_en1 = 1'b1;
				count_en2 = 1'b1;
				WE = 1'b1;
			end
			FIX: begin
				sync_clr = 1'b1;
			end
		endcase
	end
endmodule

// $Id: $
// File name:   s_box_lookup.sv
// Created:     4/11/2017
// Author:      Gabriel Chen
// Lab Section: 337-03
// Version:     1.0  Initial Design Entry
// Description: Module for the s-box lookup table
module s_box_lookup
(
  input wire [7:0] input_word,
  output reg [7:0] substituted_word
);

always_comb begin :SBOX

  case(input_word)

	0 : substituted_word = 99;
	1 : substituted_word = 124;
	2 : substituted_word = 119;
	3 : substituted_word = 123;
	4 : substituted_word = 242;
	5 : substituted_word = 107;
	6 : substituted_word = 111;
	7 : substituted_word = 197;
	8 : substituted_word = 48;
	9 : substituted_word = 1;
	10 : substituted_word = 103;
	11 : substituted_word = 43;
	12 : substituted_word = 254;
	13 : substituted_word = 215;
	14 : substituted_word = 171;
	15 : substituted_word = 118;
	16 : substituted_word = 202;
	17 : substituted_word = 130;
	18 : substituted_word = 201;
	19 : substituted_word = 125;
	20 : substituted_word = 250;
	21 : substituted_word = 89;
	22 : substituted_word = 71;
	23 : substituted_word = 240;
	24 : substituted_word = 173;
	25 : substituted_word = 212;
	26 : substituted_word = 162;
	27 : substituted_word = 175;
	28 : substituted_word = 156;
	29 : substituted_word = 164;
	30 : substituted_word = 114;
	31 : substituted_word = 192;
	32 : substituted_word = 183;
	33 : substituted_word = 253;
	34 : substituted_word = 147;
	35 : substituted_word = 38;
	36 : substituted_word = 54;
	37 : substituted_word = 63;
	38 : substituted_word = 247;
	39 : substituted_word = 204;
	40 : substituted_word = 52;
	41 : substituted_word = 165;
	42 : substituted_word = 229;
	43 : substituted_word = 241;
	44 : substituted_word = 113;
	45 : substituted_word = 216;
	46 : substituted_word = 49;
	47 : substituted_word = 21;
	48 : substituted_word = 4;
	49 : substituted_word = 199;
	50 : substituted_word = 35;
	51 : substituted_word = 195;
	52 : substituted_word = 24;
	53 : substituted_word = 150;
	54 : substituted_word = 5;
	55 : substituted_word = 154;
	56 : substituted_word = 7;
	57 : substituted_word = 18;
	58 : substituted_word = 128;
	59 : substituted_word = 226;
	60 : substituted_word = 235;
	61 : substituted_word = 39;
	62 : substituted_word = 178;
	63 : substituted_word = 117;
	64 : substituted_word = 9;
	65 : substituted_word = 131;
	66 : substituted_word = 44;
	67 : substituted_word = 26;
	68 : substituted_word = 27;
	69 : substituted_word = 110;
	70 : substituted_word = 90;
	71 : substituted_word = 160;
	72 : substituted_word = 82;
	73 : substituted_word = 59;
	74 : substituted_word = 214;
	75 : substituted_word = 179;
	76 : substituted_word = 41;
	77 : substituted_word = 227;
	78 : substituted_word = 47;
	79 : substituted_word = 132;
	80 : substituted_word = 83;
	81 : substituted_word = 209;
	82 : substituted_word = 0;
	83 : substituted_word = 237;
	84 : substituted_word = 32;
	85 : substituted_word = 252;
	86 : substituted_word = 177;
	87 : substituted_word = 91;
	88 : substituted_word = 106;
	89 : substituted_word = 203;
	90 : substituted_word = 190;
	91 : substituted_word = 57;
	92 : substituted_word = 74;
	93 : substituted_word = 76;
	94 : substituted_word = 88;
	95 : substituted_word = 207;
	96 : substituted_word = 208;
	97 : substituted_word = 239;
	98 : substituted_word = 170;
	99 : substituted_word = 251;
	100 : substituted_word = 67;
	101 : substituted_word = 77;
	102 : substituted_word = 51;
	103 : substituted_word = 133;
	104 : substituted_word = 69;
	105 : substituted_word = 249;
	106 : substituted_word = 2;
	107 : substituted_word = 127;
	108 : substituted_word = 80;
	109 : substituted_word = 60;
	110 : substituted_word = 159;
	111 : substituted_word = 168;
	112 : substituted_word = 81;
	113 : substituted_word = 163;
	114 : substituted_word = 64;
	115 : substituted_word = 143;
	116 : substituted_word = 146;
	117 : substituted_word = 157;
	118 : substituted_word = 56;
	119 : substituted_word = 245;
	120 : substituted_word = 188;
	121 : substituted_word = 182;
	122 : substituted_word = 218;
	123 : substituted_word = 33;
	124 : substituted_word = 16;
	125 : substituted_word = 255;
	126 : substituted_word = 243;
	127 : substituted_word = 210;
	128 : substituted_word = 205;
	129 : substituted_word = 12;
	130 : substituted_word = 19;
	131 : substituted_word = 236;
	132 : substituted_word = 95;
	133 : substituted_word = 151;
	134 : substituted_word = 68;
	135 : substituted_word = 23;
	136 : substituted_word = 196;
	137 : substituted_word = 167;
	138 : substituted_word = 126;
	139 : substituted_word = 61;
	140 : substituted_word = 100;
	141 : substituted_word = 93;
	142 : substituted_word = 25;
	143 : substituted_word = 115;
	144 : substituted_word = 96;
	145 : substituted_word = 129;
	146 : substituted_word = 79;
	147 : substituted_word = 220;
	148 : substituted_word = 34;
	149 : substituted_word = 42;
	150 : substituted_word = 144;
	151 : substituted_word = 136;
	152 : substituted_word = 70;
	153 : substituted_word = 238;
	154 : substituted_word = 184;
	155 : substituted_word = 20;
	156 : substituted_word = 222;
	157 : substituted_word = 94;
	158 : substituted_word = 11;
	159 : substituted_word = 219;
	160 : substituted_word = 224;
	161 : substituted_word = 50;
	162 : substituted_word = 58;
	163 : substituted_word = 10;
	164 : substituted_word = 73;
	165 : substituted_word = 6;
	166 : substituted_word = 36;
	167 : substituted_word = 92;
	168 : substituted_word = 194;
	169 : substituted_word = 211;
	170 : substituted_word = 172;
	171 : substituted_word = 98;
	172 : substituted_word = 145;
	173 : substituted_word = 149;
	174 : substituted_word = 228;
	175 : substituted_word = 121;
	176 : substituted_word = 231;
	177 : substituted_word = 200;
	178 : substituted_word = 55;
	179 : substituted_word = 109;
	180 : substituted_word = 141;
	181 : substituted_word = 213;
	182 : substituted_word = 78;
	183 : substituted_word = 169;
	184 : substituted_word = 108;
	185 : substituted_word = 86;
	186 : substituted_word = 244;
	187 : substituted_word = 234;
	188 : substituted_word = 101;
	189 : substituted_word = 122;
	190 : substituted_word = 174;
	191 : substituted_word = 8;
	192 : substituted_word = 186;
	193 : substituted_word = 120;
	194 : substituted_word = 37;
	195 : substituted_word = 46;
	196 : substituted_word = 28;
	197 : substituted_word = 166;
	198 : substituted_word = 180;
	199 : substituted_word = 198;
	200 : substituted_word = 232;
	201 : substituted_word = 221;
	202 : substituted_word = 116;
	203 : substituted_word = 31;
	204 : substituted_word = 75;
	205 : substituted_word = 189;
	206 : substituted_word = 139;
	207 : substituted_word = 138;
	208 : substituted_word = 112;
	209 : substituted_word = 62;
	210 : substituted_word = 181;
	211 : substituted_word = 102;
	212 : substituted_word = 72;
	213 : substituted_word = 3;
	214 : substituted_word = 246;
	215 : substituted_word = 14;
	216 : substituted_word = 97;
	217 : substituted_word = 53;
	218 : substituted_word = 87;
	219 : substituted_word = 185;
	220 : substituted_word = 134;
	221 : substituted_word = 193;
	222 : substituted_word = 29;
	223 : substituted_word = 158;
	224 : substituted_word = 225;
	225 : substituted_word = 248;
	226 : substituted_word = 152;
	227 : substituted_word = 17;
	228 : substituted_word = 105;
	229 : substituted_word = 217;
	230 : substituted_word = 142;
	231 : substituted_word = 148;
	232 : substituted_word = 155;
	233 : substituted_word = 30;
	234 : substituted_word = 135;
	235 : substituted_word = 233;
	236 : substituted_word = 206;
	237 : substituted_word = 85;
	238 : substituted_word = 40;
	239 : substituted_word = 223;
	240 : substituted_word = 140;
	241 : substituted_word = 161;
	242 : substituted_word = 137;
	243 : substituted_word = 13;
	244 : substituted_word = 191;
	245 : substituted_word = 230;
	246 : substituted_word = 66;
	247 : substituted_word = 104;
	248 : substituted_word = 65;
	249 : substituted_word = 153;
	250 : substituted_word = 45;
	251 : substituted_word = 15;
	252 : substituted_word = 176;
	253 : substituted_word = 84;
	254 : substituted_word = 187;
	255 : substituted_word = 22;

  endcase
end

endmodule


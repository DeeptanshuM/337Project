// $Id: $
// File name:   tb_rcv_fifo.sv
// Created:     4/15/2017
// Author:      Natat Sombuntham
// Lab Section: 337-03
// Version:     1.0  Initial Design Entry
// Description: Test bench for top level module rcv_fifo/
`timescale 1ns / 10ps
module tb_rcv_fifo();
	parameter CLK_PERIOD				= 4;
	
	reg tb_clk;
	reg tb_n_rst;
	reg [31:0] tb_HWDATA;
	reg tb_rcv_deq;
	reg tb_rcv_enq_word;
	reg tb_fix_error;
	reg [127:0] tb_rcv_fifo_out;
	reg tb_full;
	reg tb_empty;
	reg tb_framing_error;

	integer tb_test_case_num;

	rcv_fifo DUT
	(
		.clk(tb_clk),
		.n_rst(tb_n_rst),
		.HWDATA(tb_HWDATA),
		.rcv_deq(tb_rcv_deq),
		.rcv_enq_word(tb_rcv_enq_word),
		.fix_error(tb_fix_error),
		.rcv_fifo_out(tb_rcv_fifo_out),
		.full(tb_full),
		.empty(tb_empty),
		.framing_error(tb_framing_error)
	);

	always
	begin : CLK_GEN
		tb_clk = 1'b0;
		#(CLK_PERIOD / 2.0);
		tb_clk = 1'b1;
		#(CLK_PERIOD / 2.0);
	end

	task reset_dut;
	begin
		// Activate the design's reset (does not need to be synchronize with clock)
		tb_n_rst = 1'b0;
		
		// Wait for a couple clock cycles
		@(posedge tb_clk);
		@(posedge tb_clk);
		
		// Release the reset
		@(negedge tb_clk);
		tb_n_rst = 1'b1;
		
		// Wait for a while before activating the design
		@(posedge tb_clk);
		@(posedge tb_clk);
	end
	endtask

	task chk_full_empty_error;
		input exp_full;
		input exp_empty;
		input exp_error;
	begin
		assert(exp_full == tb_full)
		begin
			$info("Test Case #%0d: Had a correct FIFO FULL value", tb_test_case_num);
		end else begin
			$error("Test Case #%0d: Had an incorrect FIFO FULL value ******************************", tb_test_case_num);
		end
		assert(exp_empty == tb_empty)
		begin
			$info("Test Case #%0d: Had a correct FIFO EMPTY value", tb_test_case_num);
		end else begin
			$error("Test Case #%0d: Had an incorrect FIFO EMPTY value ******************************", tb_test_case_num);
		end
		assert(exp_error == tb_framing_error)
		begin
			$info("Test Case #%0d: Had a correct FIFO ERROR value", tb_test_case_num);
		end else begin
			$error("Test Case #%0d: Had an incorrect FIFO ERROR value ******************************", tb_test_case_num);
		end
	end
	endtask

	task send_data;
		input [31:0] data;
	begin
		@(negedge tb_clk);
		tb_HWDATA = data;
		tb_rcv_enq_word = 1'b1;
		@(negedge tb_clk);
		tb_rcv_enq_word = 1'b0;
	end
	endtask

	task send_burst;
		input [127:0] data;
	begin
		@(negedge tb_clk);
		tb_rcv_enq_word = 1'b1;
		tb_HWDATA = data[127:96];
		@(negedge tb_clk);
		tb_HWDATA = data[95:64];
		@(negedge tb_clk);
		tb_HWDATA = data[63:32];
		@(negedge tb_clk);
		tb_HWDATA = data[31:0];
		@(negedge tb_clk);
		tb_rcv_enq_word = 1'b0;
		@(negedge tb_clk);

	end
	endtask
	task send_burst_all;
		input [127:0] data1;
		input [127:0] data2;
		input [127:0] data3;
	begin
		@(negedge tb_clk);
		tb_rcv_enq_word = 1'b1;
		tb_HWDATA = data1[127:96];
		@(negedge tb_clk);
		tb_HWDATA = data1[95:64];
		@(negedge tb_clk);
		tb_HWDATA = data1[63:32];
		@(negedge tb_clk);
		tb_HWDATA = data1[31:0];
		@(negedge tb_clk);
		tb_HWDATA = data2[127:96];
		@(negedge tb_clk);
		tb_HWDATA = data2[95:64];
		@(negedge tb_clk);
		tb_HWDATA = data2[63:32];
		@(negedge tb_clk);
		tb_HWDATA = data2[31:0];
		@(negedge tb_clk);
		tb_HWDATA = data3[127:96];
		@(negedge tb_clk);
		tb_HWDATA = data3[95:64];
		@(negedge tb_clk);
		tb_HWDATA = data3[63:32];
		@(negedge tb_clk);
		tb_HWDATA = data3[31:0];
		@(negedge tb_clk);
		tb_rcv_enq_word = 1'b0;
		@(negedge tb_clk);

	end
	endtask

	task deq_data;
	begin
		@(negedge tb_clk);
		tb_rcv_deq = 1'b1;
		@(negedge tb_clk);
		tb_rcv_deq = 1'b0;
		@(negedge tb_clk);
	end
	endtask

	task deq_burst;
	begin
		@(negedge tb_clk);
		tb_rcv_deq = 1'b1;
		@(negedge tb_clk);
		@(negedge tb_clk);
		@(negedge tb_clk);
		tb_rcv_deq = 1'b0;
		@(negedge tb_clk);
	end
	endtask

	task chk_output;
		input [127:0] data;
	begin
		assert(data == tb_rcv_fifo_out)
		begin
			$info("Test Case #%0d: Had a correct FIFO DATA value", tb_test_case_num);
		end else begin
			$error("Test Case #%0d: Had an incorrect FIFO DATA value ******************************", tb_test_case_num);
		end
	end
	endtask
	
	reg e_full;
	reg e_empty;
	reg e_error;
	initial begin
		tb_rcv_deq = 1'b0;
		tb_rcv_enq_word = 1'b0;
		tb_fix_error = 1'b0;		
		tb_n_rst = 1'b1;
		tb_test_case_num = 0;
		//TEST 0 TEST AFTER RESET
		reset_dut();
		e_full = 1'b0;
		e_empty = 1'b1;
		e_error = 1'b0;
		chk_full_empty_error(e_full, e_empty, e_error);
		tb_test_case_num = tb_test_case_num + 1;


		//TEST1 TEST AFTER ONE ENQUEUE
		send_data(32'hAA);
		e_full = 1'b0;
		e_empty = 1'b0;
		e_error = 1'b1;
		@(negedge tb_clk);
		chk_full_empty_error(e_full, e_empty, e_error);
		tb_test_case_num = tb_test_case_num + 1;

		//TEST2 TEST AFTER THREE MORE ENQUEUES
		send_data(32'hBB);
		send_data(32'hCC);
		send_data(32'hDD);
		e_full = 1'b0;
		e_empty = 1'b0;
		e_error = 1'b0;
		@(negedge tb_clk);
		chk_full_empty_error(e_full, e_empty, e_error);
		chk_output({32'hAA, 32'hBB, 32'hCC, 32'hDD});
		tb_test_case_num = tb_test_case_num + 1;

		//TEST3 TEST AFTER ONE DEQUEUE
		deq_data();
		e_full = 1'b0;
		e_empty = 1'b1;
		e_error = 1'b0;
		@(negedge tb_clk);
		chk_full_empty_error(e_full, e_empty, e_error);
		tb_test_case_num = tb_test_case_num + 1;

		//TEST4 TEST AFTER SENDING BURST
		send_burst({32'h11, 32'h22, 32'h33, 32'h44});
		chk_output({32'h11, 32'h22, 32'h33, 32'h44});
		e_full = 1'b0;
		e_empty = 1'b0;
		e_error = 1'b0;
		@(negedge tb_clk);
		chk_full_empty_error(e_full, e_empty, e_error);
		tb_test_case_num = tb_test_case_num + 1;


		//TEST5 TEST deq
		deq_data();
		e_full = 1'b0;
		e_empty = 1'b1;
		e_error = 1'b0;
		@(negedge tb_clk);
		chk_full_empty_error(e_full, e_empty, e_error);
		tb_test_case_num = tb_test_case_num + 1;

		//TEST4 TEST AFTER SENDING BURST
		send_burst_all({32'h11, 32'h22, 32'h33, 32'h44},
			       {32'h55, 32'h66, 32'h77, 32'h88},
			       {32'h99, 32'hAA, 32'hBB, 32'hCC});
		chk_output({32'h11, 32'h22, 32'h33, 32'h44});
		e_full = 1'b1;
		e_empty = 1'b0;
		e_error = 1'b0;
		@(negedge tb_clk);
		chk_full_empty_error(e_full, e_empty, e_error);
		tb_test_case_num = tb_test_case_num + 1;

		//TEST5 DEQ BURST
		deq_burst();
		e_full = 1'b0;
		e_empty = 1'b1;
		e_error = 1'b0;
		@(negedge tb_clk);
		chk_full_empty_error(e_full, e_empty, e_error);


		//TEST4 TEST AFTER SENDING BURST
		send_burst_all("A",
			       "B",
			       "C");
		e_full = 1'b1;
		e_empty = 1'b0;
		e_error = 1'b0;
		@(negedge tb_clk);
		chk_full_empty_error(e_full, e_empty, e_error);
		deq_burst();
		tb_test_case_num = tb_test_case_num + 1;
	end
	
endmodule

module byte_sub
  (
   input [127:0] lu_table,
   input [7:0] data_i,
   output [7:0]	 data_o
   );

   always_comb begin : MULTIPLEXER
      case(data_i)
	
      endcase
     end

   
     
endmodule

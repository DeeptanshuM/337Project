mg85@ecegrid-thin1.ecn.purdue.edu.3835:1489747261
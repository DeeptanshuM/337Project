// $Id: $
// File name:   tb_aes_block.sv
// Created:     4/15/2017
// Author:      Kent Gauen
// Lab Section: 337-03
// Version:     1.0  Initial Design Entry
// Description: Test bench for top level module aes_block/
`timescale 1ns / 10ps
module tb_aes_block();
	parameter CLK_PERIOD				= 4;
	
	initial begin
	   #(CLK_PERIOD);
	   
	end
	
endmodule

// AES: mix columns 

module mix_columns
  (
   input wire 	       i_mode,
   input wire [127:0]  i_data,
   output wire [127:0] o_data
   );
   
   // NOT IMPLEMENTED
   assign o_data = i_data;
   

endmodule

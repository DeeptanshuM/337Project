// $Id: $
// File name:   ahb_regs.sv
// Created:     4/18/2017
// Author:      Natat Sombuntham
// Lab Section: 337-03
// Version:     1.0  Initial Design Entry
// Description: Place to store the registers as outputs of AHB.
module ahb_regs (
	input wire       HCLK,
	input wire       HRESETn,
	input wire          HSELx,
	input wire  [31:0]  HADDR,
	input wire  [ 2:0]  HBURST,
	input wire  [ 3:0]  HPROT,
	input wire  [ 2:0]  HSIZE,
	input wire  [ 1:0]  HTRANS,
	input wire          HWRITE,
	input wire 	 key_done,
	input wire       rcv_fifo_full,
	input wire       rcv_fifo_empty,
	input wire       tx_fifo_empty,
	output reg       rcv_enq_word,
	output reg       tx_deq_word,
	output reg       is_encrypt_pulse,
	output reg       is_decrypt_pulse,
	output reg       key_in,
	output reg       is_status,
	output reg       HREADY,
	output reg [1:0] HRESP
);
	parameter SINGLE = 3'b000;
	parameter INCR = 3'b001;
	parameter BUZ = 2'b01;
	parameter NONSEQ = 2'b10;
	parameter SEQ = 2'b11;
	typedef enum bit [3:0] {NOP, OUTPUT_BUR, INPUT_BUR, KEY_BUR, LAST_KEY_WORD_BUR, GET_STATUS,
				ENCRYPT, DECRYPT, BUSY, ERROR, OUTPUT_BUR_BUSY, INPUT_BUR_BUSY, KEY_BUR_BUSY} opcodeType;
	typedef enum bit [2:0] {IDLE, ERR1, ERR2, BEEZ, OUT_BUR_BUSY, IN_BUR_BUSY, K_BUR_BUSY} errType;

	errType state;
	errType nextState;

//	reg tmp_rcv_enq_word;
//	reg tmp_tx_deq_word;
	reg tmp_is_encrypt_pulse;
	reg tmp_is_decrypt_pulse;
	reg tmp_key_in;
	reg tmp_is_status;
	reg [ 3:0]  opcode;
	
	always_ff @ (negedge HRESETn, posedge HCLK) begin 
		if (HRESETn == 1'b0) begin
			is_encrypt_pulse <= 1'b0;
			is_decrypt_pulse <= 1'b0;
			key_in <= 1'b0;
			is_status <= 1'b0;
		end else begin
			is_encrypt_pulse <= tmp_is_encrypt_pulse;
			is_decrypt_pulse <= tmp_is_decrypt_pulse;
			key_in <= tmp_key_in;
			is_status <= tmp_is_status;
		end
	end

	always_ff @ (negedge HRESETn, posedge HCLK) begin : FSM_LOGIC
		if (HRESETn == 1'b0) begin
			state <= IDLE;
		end else begin
			state <= nextState;
		end
	end

	always_comb begin : NXT_ST_LOGIC
		nextState = state;
		case (state)
			IDLE: begin
				if (opcode == ERROR) begin
					nextState = ERR1;
				end
				else if (opcode == BUSY) begin
					nextState = BEEZ;
				end
				else if (opcode == OUTPUT_BUR_BUSY) begin
					nextState = OUT_BUR_BUSY;
				end
				else if (opcode == INPUT_BUR_BUSY) begin
					nextState = IN_BUR_BUSY;
				end
				else if (opcode == KEY_BUR_BUSY) begin
					nextState = K_BUR_BUSY;
				end
			end
			ERR1: begin
				nextState = ERR2;
			end
			ERR2: begin
				nextState = IDLE;
			end
			BEEZ: begin
				if (HTRANS != BUZ) begin
					nextState = IDLE;
				end
			end
			OUT_BUR_BUSY: begin
				if (!tx_fifo_empty) begin
					nextState = IDLE;
				end
			end
			IN_BUR_BUSY: begin
				if (!rcv_fifo_full) begin
					nextState = IDLE;
				end
			end
			K_BUR_BUSY: begin
				if (rcv_fifo_empty) begin
					nextState = IDLE;
				end
			end
		endcase
	end

	always_comb begin : OUTPUT_LOGIC
		HREADY = 1'b1;
		HRESP = 2'b00;
		case (state)
			IDLE: begin
				//do nothing
			end
			ERR1: begin
				HREADY = 1'b0;
				HRESP = 2'b01;
			end
			ERR2: begin
				HREADY = 1'b1;
				HRESP = 2'b01;
			end
			BEEZ: begin
				HREADY = 1'b0;
			end
			OUT_BUR_BUSY: begin
				HREADY = 1'b0;
			end
			IN_BUR_BUSY: begin
				HREADY = 1'b0;
			end
			K_BUR_BUSY: begin
				HREADY = 1'b0;
			end
		endcase
	end


	always_comb begin
//		tmp_rcv_enq_word = 1'b0;
		rcv_enq_word = 1'b0;
		//tmp_tx_deq_word = 1'b0;
		tx_deq_word = 1'b0;
		tmp_is_encrypt_pulse = 1'b0;
		tmp_is_decrypt_pulse = 1'b0;
		tmp_key_in = 1'b0;
		tmp_is_status = 1'b0;
		opcode = NOP;
		if (HSELx == 1'b0 || HTRANS == IDLE) begin
			//
		end
		else if (HSIZE != 2 || ((HADDR >= 32'h80 && HADDR < 32'hE0  || HADDR >= 32'h40 && HADDR < 32'h80) && key_done == 1'b0)) begin
//		else if (HSIZE != 2) begin
			opcode = ERROR;
		end
		else if (HADDR >= 32'h80 && HADDR < 32'hE0 && !HWRITE && HBURST == INCR && HTRANS != BUSY && !tx_fifo_empty) begin
			//tmp_tx_deq_word = 1'b1; //op = OUTPUT_BUR;
			tx_deq_word = 1'b1;
		end
		else if (HADDR >= 32'h80 && HADDR < 32'hE0 && !HWRITE && HBURST == INCR && HTRANS != BUSY && tx_fifo_empty) begin
			opcode = OUTPUT_BUR_BUSY;
		end
		else if (HADDR >= 32'h40 && HADDR < 32'h80 && HWRITE && HBURST == INCR && HTRANS != BUSY && !rcv_fifo_full) begin
			//tmp_rcv_enq_word = 1'b1;
			rcv_enq_word = 1'b1;// op = INPUT_BUR;
		end
		else if (HADDR >= 32'h40 && HADDR < 32'h80 && HWRITE && HBURST == INCR && HTRANS != BUSY && rcv_fifo_full) begin
			opcode = INPUT_BUR_BUSY;
		end
		else if (HADDR == 32'h10 && HWRITE && HBURST == INCR && HTRANS != BUSY && rcv_fifo_empty) begin
			//tmp_rcv_enq_word = 1'b1;  //op = KEY_BUR;
			rcv_enq_word = 1'b1;
		end
		else if (HADDR == 32'h10 && HWRITE && HBURST == INCR && HTRANS != BUSY && !rcv_fifo_empty) begin
			opcode = KEY_BUR_BUSY;
		end
		else if (HADDR >= 32'h14 && HADDR < 32'h1C && HWRITE && HBURST == INCR && HTRANS != BUSY) begin
//			tmp_rcv_enq_word = 1'b1;  //op = KEY_BUR;
			rcv_enq_word = 1'b1;
		end
		else if (HADDR == 32'h1C && HWRITE && HBURST == INCR && HTRANS != BUSY) begin
//			tmp_rcv_enq_word = 1'b1;  //op = KEY_BUR;
			rcv_enq_word = 1'b1;
			tmp_key_in = 1'b1;
			//op = LAST_KEY_WORD_BUR;
		end
		else if (HADDR == 32'h00 && !HWRITE && HBURST == SINGLE && HTRANS == NONSEQ) begin
			tmp_is_status = 1'b1;//op = GET_STATUS;
		end
		else if (HADDR == 32'h04 && HWRITE && HBURST == SINGLE && HTRANS == NONSEQ) begin
			tmp_is_encrypt_pulse = 1'b1;//op = ENCRYPT;
		end
		else if (HADDR == 32'h08 && HWRITE && HBURST == SINGLE && HTRANS == NONSEQ) begin
			tmp_is_decrypt_pulse = 1'b1; //op = DECRYPT;
		end
		else if (HTRANS == BUZ) begin
			opcode = BUSY;
		end
		else begin
			opcode = ERROR;
		end
	end
endmodule

// $Id: $
// File name:   ahb_address_decoder.sv
// Created:     4/18/2017
// Author:      Natat Sombuntham
// Lab Section: 337-03
// Version:     1.0  Initial Design Entry
// Description: Decoder for address.

module ahb_address_decoder (
	input wire          HSELx,
	input wire  [31:0]  HADDR,
	input wire  [ 2:0]  HBURST,
	input wire  [ 3:0]  HPROT,
	input wire  [ 2:0]  HSIZE,
	input wire  [ 1:0]  HTRANS,
	input wire          HWRITE,
	input wire          rcv_fifo_full,
	input wire          rcv_fifo_empty,
	input wire          tx_fifo_empty,
	output wire [ 3:0]  opcode
);
	parameter SINGLE = 3'b000;
	parameter INCR = 3'b001;
	parameter IDLE = 2'b00;
	parameter BUZ = 2'b01;
	parameter NONSEQ = 2'b10;
	parameter SEQ = 2'b11;

	typedef enum bit [3:0] {NOP, OUTPUT_BUR, INPUT_BUR, KEY_BUR, LAST_KEY_WORD_BUR, GET_STATUS,
				ENCRYPT, DECRYPT, BUSY, ERROR, OUTPUT_BUR_BUSY, INPUT_BUR_BUSY, KEY_BUR_BUSY} opcodeType;
	opcodeType op;
	assign opcode = op;
	always_comb begin
		if (HSELx == 1'b0 || HTRANS == IDLE) begin
			op = NOP;
		end
		else if (HSIZE != 2) begin
			op = ERROR;
		end
		else if (HADDR >= 32'h80 && HADDR < 32'hE0 && !HWRITE && HBURST == INCR && HTRANS != BUSY && !tx_fifo_empty) begin
			op = OUTPUT_BUR;
		end
		else if (HADDR >= 32'h80 && HADDR < 32'hE0 && !HWRITE && HBURST == INCR && HTRANS != BUSY && tx_fifo_empty) begin
			op = OUTPUT_BUR_BUSY;
		end
		else if (HADDR >= 32'h40 && HADDR < 32'h80 && HWRITE && HBURST == INCR && HTRANS != BUSY && !rcv_fifo_full) begin
			op = INPUT_BUR;
		end
		else if (HADDR >= 32'h40 && HADDR < 32'h80 && HWRITE && HBURST == INCR && HTRANS != BUSY && rcv_fifo_full) begin
			op = INPUT_BUR_BUSY;
		end
		else if (HADDR == 32'h10 && HWRITE && HBURST == INCR && HTRANS != BUSY && rcv_fifo_empty) begin
			op = KEY_BUR;
		end
		else if (HADDR == 32'h10 && HWRITE && HBURST == INCR && HTRANS != BUSY && !rcv_fifo_empty) begin
			op = KEY_BUR_BUSY;
		end
		else if (HADDR >= 32'h14 && HADDR < 32'h1C && HWRITE && HBURST == INCR && HTRANS != BUSY) begin
			op = KEY_BUR;
		end
		else if (HADDR == 32'h1C && HWRITE && HBURST == INCR && HTRANS != BUSY) begin
			op = LAST_KEY_WORD_BUR;
		end
		else if (HADDR == 32'h00 && !HWRITE && HBURST == SINGLE && HTRANS == NONSEQ) begin
			op = GET_STATUS;
		end
		else if (HADDR == 32'h04 && HWRITE && HBURST == SINGLE && HTRANS == NONSEQ) begin
			op = ENCRYPT;
		end
		else if (HADDR == 32'h08 && HWRITE && HBURST == SINGLE && HTRANS == NONSEQ) begin
			op = DECRYPT;
		end
		else if (HTRANS == BUZ) begin
			op = BUSY;
		end
		else begin
			op = ERROR;
		end
	end
endmodule
